grammar edu:umn:cs:melt:exts:ableC:regex:mda_test;

import edu:umn:cs:melt:ableC:host;

copper_mda testConcreteSyntax(ablecParser) {
  edu:umn:cs:melt:exts:ableC:regex:concreteSyntax;
}
