grammar edu:umn:cs:melt:exts:ableC:regex;

exports edu:umn:cs:melt:exts:ableC:regex:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:regex:concretesyntax;